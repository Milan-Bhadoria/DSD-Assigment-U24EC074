`timescale 1ns / 1ps
module LUT_ram #(parameter W = 32,
      D = 16384
)(
   input clk,write_en,
   input [W-1:0]data_in,
   input [$clog2(D)-1:0]write_addr,read_addr,
   output reg [W-1:0] out
);
  reg [W-1:0] lut[D-1:0];
  always@(posedge clk)begin
     if(write_en)begin
       lut[write_addr] <= data_in;
     end
   else out <= lut[read_addr];
   end
endmodule
